module vmate5

struct NullGrammar {
	Grammar
	name       string = 'Null Grammar'
	scope_name string = 'text.plain.null-grammar'
}
